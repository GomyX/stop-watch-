module STOPWATCH( input logic  MAINCLOCK,MAINPUSHR,MAINPUSHL,MAINDIP1S,MAINDIP2M,
output logic [7:0] DIGIT7SEG,
output logic [3:0] ENABLE7SEG);

wire CLOCK1sec,RESETFORERROR,MODE_COUNTER,LOAD_COUNTER,STRT_COUNTER,IS_THERE_ERROR,RESET;
wire [3:0] MCOUNT0,MCOUNT1,MCOUNT2,MCOUNT3,MERROR0,MERROR1,MERROR2,MERROR3,MAINSVNSG0,MAINSVNSG1,MAINSVNSG2,MAINSVNSG3;

clkdiv CLOCKTO1SEC(MAINPUSHR, MAINCLOCK, CLOCK1sec);

MAINFSM MYFSM (CLOCK1sec,MAINPUSHR,MAINDIP1S,MAINDIP2M,MAINPUSHL,RESETFORERROR,MODE_COUNTER,LOAD_COUNTER,STRT_COUNTER,IS_THERE_ERROR,MERROR0,MERROR1,MERROR2,MERROR3);
or rstat (RESET, RESETFORERROR,MAINPUSHR);

MIN_SEC_COUNTER MYCLKCOUNT( MODE_COUNTER,STRT_COUNTER,CLOCK,CLOCK1sec, RESET,LOAD_COUNTER, MCOUNT0,MCOUNT1,MCOUNT2,MCOUNT3);

Todisplay MYDISPLAY (IS_THERE_ERROR, MCOUNT0,MCOUNT1,MCOUNT2,MCOUNT3, MERROR0,MERROR1,MERROR2,MERROR3, MAINSVNSG0,MAINSVNSG1,MAINSVNSG2,MAINSVNSG3);

disp_hex_mux finaldisplay( MAINCLOCK, MAINPUSHR, MAINSVNSG0,MAINSVNSG1,MAINSVNSG2,MAINSVNSG3 ,4'b0000 ,DIGIT7SEG, ENABLE7SEG) ;
endmodule
